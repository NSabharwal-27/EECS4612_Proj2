//====================================
// mem_resp_inf.sv
//====================================
// requests data from MEM

module mem_resp_inf(

);


endmodule