//====================================
// mem_resp_inf.sv
//====================================
// requests data from MEM

module mem_resp_inf(
    input     logic     mem_resp_valid_i,
);


endmodule